module conv_top #(
    parameter
) (
    ports
);
    
endmodule